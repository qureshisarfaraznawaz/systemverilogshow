interface svs_if (input clk, input resetn);
   logic [31:0] bus32;
endinterface
