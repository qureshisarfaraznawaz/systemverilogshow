class classA;

   function new();
   endfunction

   function void tellme();
      $display("\n\n ***************** priviet ***************\n\n");
   endfunction

endclass : classA
