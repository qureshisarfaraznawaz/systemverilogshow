class top;

   virtual

endclass : top

